-- Laboratorio 8: Contador con reset asíncrono, enable, carga, valor máximo e indicador fin de cuenta
-- Autor: María Espinosa Astilleros
-- Desarrollo: Diseñar un contador creciente de 4 bits (Q) con reset asincrono activo a nivel bajo (resetn), señal de habilitación (en),
--             valor máximo del contador (max) que puede ser inferior a 15, señal de carga activa a nivel alto (ld) que carga el valor 
--             presente en un registro R. El contador incluirá un indicador de fin de cuenta (cout) que se activará cada vez que el 
--             contador alcance el valor de fin de cuenta. 

